module InstructionMemory(
    input logic [31:0] a,
	output logic [31:0] rd
);

  // Define the ROM array with initial values
  logic [31:0] ROM [63:0];

	 // Initialize ROM with values
	initial begin
		ROM[0] = 32'b11100000010011110000000000001111;
		ROM[1] = 32'b11100010100000000000000000000010;
		ROM[2] = 32'b11100011101000001010000000010100;
		ROM[3] = 32'b11100000010011110001000000001111;
		ROM[4] = 32'b11100001010110100000000000000001;
		ROM[5] = 32'b00001010000000000000000000000101;
		ROM[6] = 32'b11100010100000010010000000000000;
		ROM[7] = 32'b11100000000000100011000000000000;
		ROM[8] = 32'b11100111100000010011000000000000;
		ROM[9] = 32'b11100111100000010011000000000000;
		ROM[10] = 32'b11100010100000010001000000000001;
		ROM[11] = 32'b11101000000000000000000000001001;
		ROM[12] = 32'b11100010100000010001000001100100;
		for (int i = 13; i < 64; i++) begin
		  ROM[i] = 32'b0;
		end
	end
	// Assign the output based on the input address
	assign rd = ROM[a[31:2]]; // word aligned
endmodule