module InstructionMemory #(parameter WIDTH = 8)
(
    input logic [WIDTH-1:0] a,
	output logic [WIDTH-1:0] rd
);

  // Define the ROM array with initial values
  logic [WIDTH-1:0] ROM [63:0];

	 // Initialize ROM with values
	initial begin
		ROM[0] = 64'b1110001110100000000001000000000000000000000000000000000000000001;
		ROM[1] = 64'b1110001010000000100000000000000000000000000000000000000000000010;
		ROM[2] = 64'b1110001110100000001010000000000000000000000000000000000000010100;
		ROM[3] = 64'b1110000101000101000000000000000000000000000000000000000000000001;
		ROM[4] = 64'b0000101000000000000000000000000000000000000000000000000000010100;
		ROM[5] = 64'b1110001010000000100010000000000000000000000000000000000000000000;
		ROM[6] = 64'b1110000000000001000011000000000000000000000000000000000000000000;
		ROM[7] = 64'b1110010000000000100011000000000000000000000000000000000000000000;
		ROM[8] = 64'b1110011000000000100100000000000000000000000000000000000000000000;
		ROM[9] = 64'b1110001010000000100001000000000000000000000000000000000000000001;
		ROM[10] = 64'b1110100000000000000000000000000000000000000000000000000000100100;
		ROM[11] = 64'b1110001010000000100001000000000000000000000000000000000001100100;
		ROM[12] = 64'b1110001010000000100001000000000000000000000000000000000001100100;
		for (int i = 13; i < 64; i++) begin
		  ROM[i] = 64'b0;
		end
	end
	// Assign the output based on the input address
	assign rd = ROM[a[63:2]]; // word aligned
endmodule